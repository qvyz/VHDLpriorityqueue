library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.MATH_REAL.all;


package sorter_pkg is
    type outarray is array(natural range<>) of integer;
    constant constval : integer := 11;
end package;